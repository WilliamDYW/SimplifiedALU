`timescale 1ns/1ps

module alu_test;

reg[31:0] i_datain,gr1,gr2;

wire [31:0] c;
wire zero;
wire overflow;
wire neg;

alu testalu(i_datain,gr1,gr2,c,branch,load,store);

initial
begin

$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  :zero:overflow:neg:branch:load:store:   hi   :   lo   ");
$monitor("   %h:%h: %h :%h:%h:%h:%h:%h:%h:  %h :    %h   : %h :   %h  :  %h :  %h  :%h:%h",
i_datain, testalu.opcode, testalu.func, gr1 , gr2, c, testalu.reg_A, testalu.reg_B, testalu.reg_C,
testalu.zf, testalu.vf, testalu.nf, testalu.branch, testalu.load, testalu.store,testalu.hi,testalu.lo);

//// logical left shift

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0000;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_1000_0000;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0000;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0001_0000_0000;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

//// logical right shift

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0010;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_1000_0010;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0010;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0001_0000_0010;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

//// arithmetic right shift

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0011;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_1000_0011;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0011;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0001_0000_0011;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

//// sllv

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;


#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
////srlv

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
////srav

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
////mult

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1000;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1000;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1000;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1010;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1000;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
////multu

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1001;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1001;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1001;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1001;

gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
////div

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1010;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1010;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1010;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1010;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
////divu

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1011;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1011;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1011;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1011;

gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

////add

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
gr1<=32'h8000_0000;
gr2<=32'hffff_0000;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
gr1<=32'h0000_0001;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
gr1<=32'h7fff_ffff;
gr2<=32'h7fff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
gr1<=32'h0000_0001;
gr2<=32'h7fff_fffe;

////addu

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
gr1<=32'h8000_0000;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
gr1<=32'h0000_0001;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
gr1<=32'h7fff_ffff;
gr2<=32'h7fff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
gr1<=32'h0000_0001;
gr2<=32'h7fff_fffe;

////sub

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
gr1<=32'h0000_0001;
gr2<=32'h0000_0001;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
gr1<=32'h0000_0002;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
gr1<=32'h7fff_ffff;
gr2<=32'h8fff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
gr1<=32'hffff_fffc;
gr2<=32'h7fff_fffe;

////subu

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
gr1<=32'h0000_0001;
gr2<=32'h0000_0001;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
gr1<=32'h0000_0002;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
gr1<=32'h7fff_ffff;
gr2<=32'h8fff_fffe;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
gr1<=32'hffff_fffc;
gr2<=32'h7fff_fffe;

////and

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0100;
gr1<=32'b0001_0010_0011_0100_1001_1010_1011_1100;
gr2<=32'b0101_0110_0111_1000_1101_1110_1111_0000;

////or

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0101;
gr1<=32'b0001_0010_0011_0100_1001_1010_1011_1100;
gr2<=32'b0101_0110_0111_1000_1101_1110_1111_0000;

////xor

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0110;
gr1<=32'b0001_0010_0011_0100_1001_1010_1011_1100;
gr2<=32'b0101_0110_0111_1000_1101_1110_1111_0000;


////nor

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0111;
gr1<=32'b0001_0010_0011_0100_1001_1010_1011_1100;
gr2<=32'b0101_0110_0111_1000_1101_1110_1111_0000;


////slt

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;

gr1<=32'hffff_fffe;
gr2<=32'hffff_ffff;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;

gr1<=32'h0000_0001;
gr2<=32'hffff_ffff;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;

gr1<=32'h0000_0001;
gr2<=32'h0000_1000;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;

gr1<=32'hffff_ffff;
gr2<=32'h0000_0001;

////sltu

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;

gr1<=32'hffff_fffe;
gr2<=32'hffff_ffff;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;

gr1<=32'h0001_0000;
gr2<=32'hffff_ffff;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;

gr1<=32'h0000_0001;
gr2<=32'h0000_1000;

#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;

gr1<=32'hffff_ffff;
gr2<=32'h0000_0001;

////beq

#10 i_datain<=32'b0001_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0001_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;
gr2<=32'hffff_ffff;

#10 i_datain<=32'b0001_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;
gr2<=32'h0000_0000;

#10 i_datain<=32'b0001_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;
gr2<=32'h0000_0001;

////bne

#10 i_datain<=32'b0001_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;
gr2<=32'hffff_fffe;

#10 i_datain<=32'b0001_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;
gr2<=32'hffff_ffff;

#10 i_datain<=32'b0001_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;
gr2<=32'h0000_0000;

#10 i_datain<=32'b0001_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;
gr2<=32'h0000_0001;

////addi

#10 i_datain<=32'b0010_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'h7fff_fffe;

#10 i_datain<=32'b0010_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;

#10 i_datain<=32'b0010_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0000;

#10 i_datain<=32'b0010_0000_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;

////addiu

#10 i_datain<=32'b0010_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'h7fff_fffe;

#10 i_datain<=32'b0010_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;

#10 i_datain<=32'b0010_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0000;

#10 i_datain<=32'b0010_0100_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;

////slti

#10 i_datain<=32'b0010_1000_0010_0010_0111_1111_1111_1111;

gr1<=32'h0000_0ffe;

#10 i_datain<=32'b0010_1000_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;

#10 i_datain<=32'b0010_1000_0010_0010_1111_1111_1111_1100;

gr1<=32'h0000_ffff;

#10 i_datain<=32'b0010_1000_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;

////sltiu

#10 i_datain<=32'b0010_1100_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_fffe;

#10 i_datain<=32'b0010_1100_0010_0010_1111_1111_1111_1111;

gr1<=32'hffff_ffff;

#10 i_datain<=32'b0010_1100_0010_0010_1111_1111_1111_1100;

gr1<=32'h0000_ffff;

#10 i_datain<=32'b0010_1100_0010_0010_1111_1111_1111_1111;

gr1<=32'h0000_0001;

////andi

#10 i_datain<=32'b0011_0000_0010_0010_1001_1010_1011_1100;
gr1<=32'b0101_0110_0111_1000_1101_1110_1111_0000;

////ori

#10 i_datain<=32'b0011_0100_0010_0010_1001_1010_1011_1100;
gr1<=32'b0101_0110_0111_1000_1101_1110_1111_0000;

////xori

#10 i_datain<=32'b0011_1000_0010_0010_1001_1010_1011_1100;
gr1<=32'b0101_0110_0111_1000_1101_1110_1111_0000;

////lw

#10 i_datain<=32'b1000_1100_0010_0010_0000_0000_0000_0001;

gr1<=32'h0800_0008;

////sw

#10 i_datain<=32'b1010_1100_0010_0010_0000_0000_0000_0001;

gr1<=32'h0800_0008;

#10 $finish;
end
endmodule